`include "riscv_no_csr_asm_program_gen.sv"