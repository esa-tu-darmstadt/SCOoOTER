package Types;
 
typedef 32 XLEN;
typedef 32 ILEN;
typedef 4 IFUINST;
typedef 2 ISSUEWIDTH;

typedef 4 RESETVEC;
typedef 'h10000 BRAMSIZE;

typedef Bit#(5) RADDR;

endpackage