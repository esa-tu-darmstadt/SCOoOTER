package Types;
 
typedef 32 XLEN;
typedef 32 ILEN;
typedef 4 IFUINST;
typedef 1 ISSUEWIDTH;

typedef 0 RESETVEC;
typedef 'h10000 BRAMSIZE;

typedef Bit#(5) RADDR;

typedef 16 ROBDEPTH;

typedef 16 INST_WINDOW;

typedef 4 NUM_FU;
typedef 4 NUM_RS;

endpackage