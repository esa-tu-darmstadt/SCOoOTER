package Fetch;

import BlueAXI :: *;
import Types :: *;
import Interfaces :: *;
import GetPut :: *;
import Inst_Types :: *;
import Decode :: *;
import FIFO :: *;
import FIFOF :: *;
import SpecialFIFOs :: *;
import MIMO :: *;
import Vector :: *;
import Debug::*;

(* synthesize *)
module mkFetch(FetchIFC) provisos(
        Mul#(XLEN, IFUINST, ifuwidth) //the width of the IFU axi must be as large as the size of a word times the issuewidth
);

    //AXI for mem access
    AXI4_Master_Rd#(XLEN, ifuwidth, 0, 0) axi <- mkAXI4_Master_Rd(0, 0, False);

    //pc points to next instruction to load
    //pc is a CREG, port 2 is used for fetching the next instruction
    // port 1 is used to redirect the program counter
    //port 0 is used to advance the PC
    Reg#(Bit#(XLEN)) pc[3] <- mkCReg(3, fromInteger(valueof(RESETVEC)));
    Reg#(UInt#(XLEN)) epoch[2] <- mkCReg(2, 0);
    FIFO#(Bit#(XLEN)) inflight_pcs <- mkPipelineFIFO();
    FIFO#(UInt#(XLEN)) inflight_epoch <- mkPipelineFIFO();
    //holds outbound Instruction and PC
    FIFOF#(Vector#(IFUINST, Tuple3#(Bit#(32), Bit#(32), UInt#(32)))) fetched_inst <- mkPipelineFIFOF();
    FIFOF#(MIMO::LUInt#(IFUINST)) fetched_amount <- mkPipelineFIFOF();


    //Requests data from memory
    //Explicit condition: Fires if the previous read has been evaluated
    // Due to the PC FIFO
    rule requestRead;
        axi4_read_data(axi, pc[2], 0);
        inflight_pcs.enq(pc[2]);
        inflight_epoch.enq(epoch[1]);
    endrule

    rule dropReadResp (inflight_epoch.first() != epoch[1]);
        let r <- axi.response.get;
        inflight_pcs.deq();
        inflight_epoch.deq();
        dbg_print(Fetch, $format("drop read"));
    endrule

    // Evaluates fetched instructions if there is enough space in the instruction window
    // TODO: make enqueued value dynamic
    rule getReadResp (inflight_epoch.first() == epoch[1]);
        let r <- axi.response.get;
        Bit#(ifuwidth) dat = r.data;
        let acqpc = inflight_pcs.first(); inflight_pcs.deq();
        inflight_epoch.deq();

        Vector#(IFUINST, Tuple3#(Bit#(32), Bit#(32), UInt#(XLEN))) instructions_v = newVector; // temporary inst storage
        
        Bit#(XLEN) startpoint = (acqpc>>2)%fromInteger(valueOf(IFUINST))*32; // pos of first useful instruction

        MIMO::LUInt#(IFUINST) amount = unpack(truncate( fromInteger(valueOf(IFUINST)) - (acqpc>>2)%fromInteger(valueOf(IFUINST)))); // how many inst were usefully extracted // TODO: make type smaller

        // Extract instructions
        // two conditions needed to keep static elaboration working
        for(Integer i = 0; i < valueOf(IFUINST); i=i+1) begin
            if(fromInteger(i) < amount) begin
                Bit#(XLEN) iword = dat[startpoint+fromInteger(i)*32+31 : startpoint+fromInteger(i)*32];
                instructions_v[i] = tuple3(iword, acqpc + (fromInteger(i)*4), inflight_epoch.first());
            end
        end

        // enq gathered instructions
        fetched_inst.enq(instructions_v);
        fetched_amount.enq(amount);

        // advance program counter
        // TODO: branch predictor
        pc[0] <= acqpc + (pack(extend(amount)) << 2);
    endrule

    function FetchedInstruction build_fetch_resp(Tuple3#(Bit#(32), Bit#(32), UInt#(XLEN)) in)
        = FetchedInstruction {instruction: tpl_1(in), pc: tpl_2(in), epoch: tpl_3(in)};

    interface imem_axi = axi.fab;

    method Action redirect(Bit#(XLEN) newpc);
        pc[1] <= newpc;
        dbg_print(Fetch, $format("Redirected: ", newpc));
        epoch[0] <= epoch[0]+1;

    endmethod
    
    interface GetS instructions;
        method FetchResponse first();
            let inst_vector = fetched_inst.first();
            let fetched_inst = Vector::map(build_fetch_resp, inst_vector);
            return FetchResponse {count: fetched_amount.first(), instructions: fetched_inst};
        endmethod
        method Action deq();
            fetched_inst.deq();
            fetched_amount.deq();
        endmethod
    endinterface


endmodule

endpackage